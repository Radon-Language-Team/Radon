module util

pub fn symlink_radon() {
	println('Symlinking...')
}