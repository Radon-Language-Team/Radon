module lexer

import structs

pub fn refine_tokens(mut app structs.App) {

	println('Got tokens to refine: ${app.all_tokens}')

}