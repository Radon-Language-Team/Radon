module main

import os
import cmd.util

fn main() {

	util.print_menu()

	if os.args.len > 1 {
		println("Under construction")
	}

}